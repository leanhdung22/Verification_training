//------------------------------------------------------------
//   Copyright 2013 Mentor Graphics Corporation
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//------------------------------------------------------------

class biquad_vseq extends uvm_sequence #(uvm_sequence_item);

`uvm_object_utils(biquad_vseq)

apb_sequencer apb;
uvm_sequencer #(signal_seq_item) signal;
biquad_reg_block rm;
biquad_env_config cfg;

// Co-efficient arrays
bit[23:0] c_a11[105];
bit[23:0] c_a12[105];
bit[23:0] c_b10[105];
bit[23:0] c_b11[105];
bit[32:0] c_b12[105];

setup_coefficients c_setup = setup_coefficients::type_id::create("c_setup");
signal_sweep_seq f_sweep = signal_sweep_seq::type_id::create("f_sweep");

function new(string name = "biquad_vseq");
  super.new(name);
endfunction

function void setup_coefficients();

  c_b10[0] = 24'h0002C1;
  c_b10[1] = 24'h000AD3;
  c_b10[2] = 24'h0029C9;
  c_b10[3] = 24'h004029;
  c_b10[4] = 24'h005ACF;
  c_b10[5] = 24'h007983;
  c_b10[6] = 24'h009C11;
  c_b10[7] = 24'h00C245;
  c_b10[8] = 24'h00EBF2;
  c_b10[9] = 24'h0118EC;
  c_b10[10] = 24'h014909;
  c_b10[11] = 24'h017C23;
  c_b10[12] = 24'h01B217;
  c_b10[13] = 24'h01EAC2;
  c_b10[14] = 24'h022605;
  c_b10[15] = 24'h0263C3;
  c_b10[16] = 24'h02A3DF;
  c_b10[17] = 24'h02E641;
  c_b10[18] = 24'h032ACF;
  c_b10[19] = 24'h049F60;
  c_b10[20] = 24'h063F81;
  c_b10[21] = 24'h080518;
  c_b10[22] = 24'h09EC35;
  c_b10[23] = 24'h0BF29E;
  c_b10[24] = 24'h0E1772;
  c_b10[25] = 24'h105AF9;
  c_b10[26] = 24'h12BE76;
  c_b10[27] = 24'h154414;
  c_b10[28] = 24'h17EEE0;
  c_b10[29] = 24'h1AC2C7;
  c_b10[30] = 24'h1DC4A1;
  c_b10[31] = 24'h20FA44;
  c_b10[32] = 24'h246A9C;
  c_b10[33] = 24'h281DC4;
  c_b10[34] = 24'h2C1D25;
  c_b10[35] = 24'h3ED371;
  c_b10[36] = 24'h3DAC66;
  c_b10[37] = 24'h3B6E69;
  c_b10[38] = 24'h3A573E;
  c_b10[39] = 24'h394524;
  c_b10[40] = 24'h3837FE;
  c_b10[41] = 24'h372FAE;
  c_b10[42] = 24'h362C17;
  c_b10[43] = 24'h352D1D;
  c_b10[44] = 24'h3432A3;
  c_b10[45] = 24'h333C8C;
  c_b10[46] = 24'h324ABE;
  c_b10[47] = 24'h315D1B;
  c_b10[48] = 24'h30738A;
  c_b10[49] = 24'h2F8DEF;
  c_b10[50] = 24'h2EAC31;
  c_b10[51] = 24'h2DCE36;
  c_b10[52] = 24'h2CF3E4;
  c_b10[53] = 24'h2C1D25;
  c_b10[54] = 24'h281DC4;
  c_b10[55] = 24'h246A9C;
  c_b10[56] = 24'h20FA44;
  c_b10[57] = 24'h1DC4A1;
  c_b10[58] = 24'h1AC2C7;
  c_b10[59] = 24'h17EEE0;
  c_b10[60] = 24'h154414;
  c_b10[61] = 24'h12BE76;
  c_b10[62] = 24'h105AF9;
  c_b10[63] = 24'h0E1772;
  c_b10[64] = 24'h0BF29E;
  c_b10[65] = 24'h09EC35;
  c_b10[66] = 24'h080518;
  c_b10[67] = 24'h063F81;
  c_b10[68] = 24'h049F60;
  c_b10[69] = 24'h032ACF;
  c_b10[70] = 24'h0129CC;
  c_b10[71] = 24'h0248C5;
  c_b10[72] = 24'h0467CC;
  c_b10[73] = 24'h056897;
  c_b10[74] = 24'h06600B;
  c_b10[75] = 24'h074E7E;
  c_b10[76] = 24'h083440;
  c_b10[77] = 24'h0911A2;
  c_b10[78] = 24'h09E6EF;
  c_b10[79] = 24'h0AB470;
  c_b10[80] = 24'h0B7A69;
  c_b10[81] = 24'h0C391D;
  c_b10[82] = 24'h0CF0CC;
  c_b10[83] = 24'h0DA1B3;
  c_b10[84] = 24'h0E4C0A;
  c_b10[85] = 24'h0EF00B;
  c_b10[86] = 24'h0F8DEA;
  c_b10[87] = 24'h1025D9;
  c_b10[88] = 24'h10B80A;
  c_b10[89] = 24'h1342DB;
  c_b10[90] = 24'h1555E2;
  c_b10[91] = 24'h1700A2;
  c_b10[92] = 24'h184F28;
  c_b10[93] = 24'h194A9A;
  c_b10[94] = 24'h19F9AC;
  c_b10[95] = 24'h1A60F1;
  c_b10[96] = 24'h1A8313;
  c_b10[97] = 24'h1A60F1;
  c_b10[98] = 24'h19F9AC;
  c_b10[99] = 24'h194A9A;
  c_b10[100] = 24'h184F28;
  c_b10[101] = 24'h1700A2;
  c_b10[102] = 24'h1555E2;
  c_b10[103] = 24'h1342DB;
  c_b10[104] = 24'h10B80A;
  c_b11[0] = 24'h000583;
  c_b11[1] = 24'h0015A6;
  c_b11[2] = 24'h005393;
  c_b11[3] = 24'h008052;
  c_b11[4] = 24'h00B59E;
  c_b11[5] = 24'h00F307;
  c_b11[6] = 24'h013822;
  c_b11[7] = 24'h01848B;
  c_b11[8] = 24'h01D7E5;
  c_b11[9] = 24'h0231D8;
  c_b11[10] = 24'h029212;
  c_b11[11] = 24'h02F847;
  c_b11[12] = 24'h03642E;
  c_b11[13] = 24'h03D585;
  c_b11[14] = 24'h044C0B;
  c_b11[15] = 24'h04C786;
  c_b11[16] = 24'h0547BF;
  c_b11[17] = 24'h05CC82;
  c_b11[18] = 24'h06559F;
  c_b11[19] = 24'h093EC0;
  c_b11[20] = 24'h0C7F03;
  c_b11[21] = 24'h100A30;
  c_b11[22] = 24'h13D86B;
  c_b11[23] = 24'h17E53C;
  c_b11[24] = 24'h1C2EE5;
  c_b11[25] = 24'h20B5F3;
  c_b11[26] = 24'h257CEC;
  c_b11[27] = 24'h2A8829;
  c_b11[28] = 24'h2FDDC1;
  c_b11[29] = 24'h35858F;
  c_b11[30] = 24'h3B8943;
  c_b11[31] = 24'h41F489;
  c_b11[32] = 24'h48D538;
  c_b11[33] = 24'h503B88;
  c_b11[34] = 24'h583A4B;
  c_b11[35] = 24'hFDA6E3;
  c_b11[36] = 24'hFB58CD;
  c_b11[37] = 24'hF6DCD3;
  c_b11[38] = 24'hF4AE7D;
  c_b11[39] = 24'hF28A49;
  c_b11[40] = 24'hF06FFC;
  c_b11[41] = 24'hEE5F5C;
  c_b11[42] = 24'hEC582E;
  c_b11[43] = 24'hEA5A3A;
  c_b11[44] = 24'hE86546;
  c_b11[45] = 24'hE67919;
  c_b11[46] = 24'hE4957C;
  c_b11[47] = 24'hE2BA37;
  c_b11[48] = 24'hE0E714;
  c_b11[49] = 24'hDF1BDF;
  c_b11[50] = 24'hDD5862;
  c_b11[51] = 24'hDB9C6C;
  c_b11[52] = 24'hD9E7C9;
  c_b11[53] = 24'hD83A4B;
  c_b11[54] = 24'hD03B88;
  c_b11[55] = 24'hC8D538;
  c_b11[56] = 24'hC1F489;
  c_b11[57] = 24'hBB8943;
  c_b11[58] = 24'hB5858F;
  c_b11[59] = 24'hAFDDC1;
  c_b11[60] = 24'hAA8829;
  c_b11[61] = 24'hA57CEC;
  c_b11[62] = 24'hA0B5F3;
  c_b11[63] = 24'h9C2EE5;
  c_b11[64] = 24'h97E53C;
  c_b11[65] = 24'h93D86B;
  c_b11[66] = 24'h900A30;
  c_b11[67] = 24'h8C7F03;
  c_b11[68] = 24'h893EC0;
  c_b11[69] = 24'h86559F;
  c_b11[70] = 24'h000000;
  c_b11[71] = 24'h000000;
  c_b11[72] = 24'h000000;
  c_b11[73] = 24'h000000;
  c_b11[74] = 24'h000000;
  c_b11[75] = 24'h000000;
  c_b11[76] = 24'h000000;
  c_b11[77] = 24'h000000;
  c_b11[78] = 24'h000000;
  c_b11[79] = 24'h000000;
  c_b11[80] = 24'h000000;
  c_b11[81] = 24'h000000;
  c_b11[82] = 24'h000000;
  c_b11[83] = 24'h000000;
  c_b11[84] = 24'h000000;
  c_b11[85] = 24'h000000;
  c_b11[86] = 24'h000000;
  c_b11[87] = 24'h000000;
  c_b11[88] = 24'h000000;
  c_b11[89] = 24'h000000;
  c_b11[90] = 24'h000000;
  c_b11[91] = 24'h000000;
  c_b11[92] = 24'h000000;
  c_b11[93] = 24'h000000;
  c_b11[94] = 24'h000000;
  c_b11[95] = 24'h000000;
  c_b11[96] = 24'h000000;
  c_b11[97] = 24'h000000;
  c_b11[98] = 24'h000000;
  c_b11[99] = 24'h000000;
  c_b11[100] = 24'h000000;
  c_b11[101] = 24'h000000;
  c_b11[102] = 24'h000000;
  c_b11[103] = 24'h000000;
  c_b11[104] = 24'h000000;
  c_b12[0] = 24'h0002C1;
  c_b12[1] = 24'h000AD3;
  c_b12[2] = 24'h0029C9;
  c_b12[3] = 24'h004029;
  c_b12[4] = 24'h005ACF;
  c_b12[5] = 24'h007983;
  c_b12[6] = 24'h009C11;
  c_b12[7] = 24'h00C245;
  c_b12[8] = 24'h00EBF2;
  c_b12[9] = 24'h0118EC;
  c_b12[10] = 24'h014909;
  c_b12[11] = 24'h017C23;
  c_b12[12] = 24'h01B217;
  c_b12[13] = 24'h01EAC2;
  c_b12[14] = 24'h022605;
  c_b12[15] = 24'h0263C3;
  c_b12[16] = 24'h02A3DF;
  c_b12[17] = 24'h02E641;
  c_b12[18] = 24'h032ACF;
  c_b12[19] = 24'h049F60;
  c_b12[20] = 24'h063F81;
  c_b12[21] = 24'h080518;
  c_b12[22] = 24'h09EC35;
  c_b12[23] = 24'h0BF29E;
  c_b12[24] = 24'h0E1772;
  c_b12[25] = 24'h105AF9;
  c_b12[26] = 24'h12BE76;
  c_b12[27] = 24'h154414;
  c_b12[28] = 24'h17EEE0;
  c_b12[29] = 24'h1AC2C7;
  c_b12[30] = 24'h1DC4A1;
  c_b12[31] = 24'h20FA44;
  c_b12[32] = 24'h246A9C;
  c_b12[33] = 24'h281DC4;
  c_b12[34] = 24'h2C1D25;
  c_b12[35] = 24'h3ED371;
  c_b12[36] = 24'h3DAC66;
  c_b12[37] = 24'h3B6E69;
  c_b12[38] = 24'h3A573E;
  c_b12[39] = 24'h394524;
  c_b12[40] = 24'h3837FE;
  c_b12[41] = 24'h372FAE;
  c_b12[42] = 24'h362C17;
  c_b12[43] = 24'h352D1D;
  c_b12[44] = 24'h3432A3;
  c_b12[45] = 24'h333C8C;
  c_b12[46] = 24'h324ABE;
  c_b12[47] = 24'h315D1B;
  c_b12[48] = 24'h30738A;
  c_b12[49] = 24'h2F8DEF;
  c_b12[50] = 24'h2EAC31;
  c_b12[51] = 24'h2DCE36;
  c_b12[52] = 24'h2CF3E4;
  c_b12[53] = 24'h2C1D25;
  c_b12[54] = 24'h281DC4;
  c_b12[55] = 24'h246A9C;
  c_b12[56] = 24'h20FA44;
  c_b12[57] = 24'h1DC4A1;
  c_b12[58] = 24'h1AC2C7;
  c_b12[59] = 24'h17EEE0;
  c_b12[60] = 24'h154414;
  c_b12[61] = 24'h12BE76;
  c_b12[62] = 24'h105AF9;
  c_b12[63] = 24'h0E1772;
  c_b12[64] = 24'h0BF29E;
  c_b12[65] = 24'h09EC35;
  c_b12[66] = 24'h080518;
  c_b12[67] = 24'h063F81;
  c_b12[68] = 24'h049F60;
  c_b12[69] = 24'h032ACF;
  c_b12[70] = 24'h8129CC;
  c_b12[71] = 24'h8248C5;
  c_b12[72] = 24'h8467CC;
  c_b12[73] = 24'h856897;
  c_b12[74] = 24'h86600B;
  c_b12[75] = 24'h874E7E;
  c_b12[76] = 24'h883440;
  c_b12[77] = 24'h8911A2;
  c_b12[78] = 24'h89E6EF;
  c_b12[79] = 24'h8AB470;
  c_b12[80] = 24'h8B7A69;
  c_b12[81] = 24'h8C391D;
  c_b12[82] = 24'h8CF0CC;
  c_b12[83] = 24'h8DA1B3;
  c_b12[84] = 24'h8E4C0A;
  c_b12[85] = 24'h8EF00B;
  c_b12[86] = 24'h8F8DEA;
  c_b12[87] = 24'h9025D9;
  c_b12[88] = 24'h90B80A;
  c_b12[89] = 24'h9342DB;
  c_b12[90] = 24'h9555E2;
  c_b12[91] = 24'h9700A2;
  c_b12[92] = 24'h984F28;
  c_b12[93] = 24'h994A9A;
  c_b12[94] = 24'h99F9AC;
  c_b12[95] = 24'h9A60F1;
  c_b12[96] = 24'h9A8313;
  c_b12[97] = 24'h9A60F1;
  c_b12[98] = 24'h99F9AC;
  c_b12[99] = 24'h994A9A;
  c_b12[100] = 24'h984F28;
  c_b12[101] = 24'h9700A2;
  c_b12[102] = 24'h9555E2;
  c_b12[103] = 24'h9342DB;
  c_b12[104] = 24'h90B80A;
  c_a11[0] = 24'hFDA160;
  c_a11[1] = 24'hFB4326;
  c_a11[2] = 24'hF68940;
  c_a11[3] = 24'hF42E2B;
  c_a11[4] = 24'hF1D4AA;
  c_a11[5] = 24'hEF7CF4;
  c_a11[6] = 24'hED2739;
  c_a11[7] = 24'hEAD3A3;
  c_a11[8] = 24'hE88255;
  c_a11[9] = 24'hE6336E;
  c_a11[10] = 24'hE3E707;
  c_a11[11] = 24'hE19D34;
  c_a11[12] = 24'hDF5608;
  c_a11[13] = 24'hDD118F;
  c_a11[14] = 24'hDACFD3;
  c_a11[15] = 24'hD890DC;
  c_a11[16] = 24'hD654AD;
  c_a11[17] = 24'hD41B47;
  c_a11[18] = 24'hD1E4AB;
  c_a11[19] = 24'hC6FCC7;
  c_a11[20] = 24'hBC5634;
  c_a11[21] = 24'hB1EA58;
  c_a11[22] = 24'hA7B0D7;
  c_a11[23] = 24'h9DA052;
  c_a11[24] = 24'h93AEDB;
  c_a11[25] = 24'h89D235;
  c_a11[26] = 24'h800000;
  c_a11[27] = 24'h09D235;
  c_a11[28] = 24'h13AEDB;
  c_a11[29] = 24'h1DA052;
  c_a11[30] = 24'h27B0D7;
  c_a11[31] = 24'h31EA58;
  c_a11[32] = 24'h3C5634;
  c_a11[33] = 24'h46FCC7;
  c_a11[34] = 24'h51E4AB;
  c_a11[35] = 24'hFDA160;
  c_a11[36] = 24'hFB4326;
  c_a11[37] = 24'hF68940;
  c_a11[38] = 24'hF42E2B;
  c_a11[39] = 24'hF1D4AA;
  c_a11[40] = 24'hEF7CF4;
  c_a11[41] = 24'hED2739;
  c_a11[42] = 24'hEAD3A3;
  c_a11[43] = 24'hE88255;
  c_a11[44] = 24'hE6336E;
  c_a11[45] = 24'hE3E707;
  c_a11[46] = 24'hE19D34;
  c_a11[47] = 24'hDF5608;
  c_a11[48] = 24'hDD118F;
  c_a11[49] = 24'hDACFD3;
  c_a11[50] = 24'hD890DC;
  c_a11[51] = 24'hD654AD;
  c_a11[52] = 24'hD41B47;
  c_a11[53] = 24'hD1E4AB;
  c_a11[54] = 24'hC6FCC7;
  c_a11[55] = 24'hBC5634;
  c_a11[56] = 24'hB1EA58;
  c_a11[57] = 24'hA7B0D7;
  c_a11[58] = 24'h9DA052;
  c_a11[59] = 24'h93AEDB;
  c_a11[60] = 24'h89D235;
  c_a11[61] = 24'h800000;
  c_a11[62] = 24'h09D235;
  c_a11[63] = 24'h13AEDB;
  c_a11[64] = 24'h1DA052;
  c_a11[65] = 24'h27B0D7;
  c_a11[66] = 24'h31EA58;
  c_a11[67] = 24'h3C5634;
  c_a11[68] = 24'h46FCC7;
  c_a11[69] = 24'h51E4AB;
  c_a11[70] = 24'hFDA160;
  c_a11[71] = 24'hFB4326;
  c_a11[72] = 24'hF68940;
  c_a11[73] = 24'hF42E2B;
  c_a11[74] = 24'hF1D4AA;
  c_a11[75] = 24'hEF7CF4;
  c_a11[76] = 24'hED2739;
  c_a11[77] = 24'hEAD3A3;
  c_a11[78] = 24'hE88255;
  c_a11[79] = 24'hE6336E;
  c_a11[80] = 24'hE3E707;
  c_a11[81] = 24'hE19D34;
  c_a11[82] = 24'hDF5608;
  c_a11[83] = 24'hDD118F;
  c_a11[84] = 24'hDACFD3;
  c_a11[85] = 24'hD890DC;
  c_a11[86] = 24'hD654AD;
  c_a11[87] = 24'hD41B47;
  c_a11[88] = 24'hD1E4AB;
  c_a11[89] = 24'hC6FCC7;
  c_a11[90] = 24'hBC5634;
  c_a11[91] = 24'hB1EA58;
  c_a11[92] = 24'hA7B0D7;
  c_a11[93] = 24'h9DA052;
  c_a11[94] = 24'h93AEDB;
  c_a11[95] = 24'h89D235;
  c_a11[96] = 24'h800000;
  c_a11[97] = 24'h09D235;
  c_a11[98] = 24'h13AEDB;
  c_a11[99] = 24'h1DA052;
  c_a11[100] = 24'h27B0D7;
  c_a11[101] = 24'h31EA58;
  c_a11[102] = 24'h3C5634;
  c_a11[103] = 24'h46FCC7;
  c_a11[104] = 24'h51E4AB;
  c_a12[0] = 24'h3DAC66;
  c_a12[1] = 24'h3B6E74;
  c_a12[2] = 24'h373067;
  c_a12[3] = 24'h352ED0;
  c_a12[4] = 24'h333FE8;
  c_a12[5] = 24'h316303;
  c_a12[6] = 24'h2F977E;
  c_a12[7] = 24'h2DDCBA;
  c_a12[8] = 24'h2C3220;
  c_a12[9] = 24'h2A971F;
  c_a12[10] = 24'h290B2C;
  c_a12[11] = 24'h278DC4;
  c_a12[12] = 24'h261E66;
  c_a12[13] = 24'h24BC99;
  c_a12[14] = 24'h2367EA;
  c_a12[15] = 24'h221FE8;
  c_a12[16] = 24'h20E42B;
  c_a12[17] = 24'h1FB44C;
  c_a12[18] = 24'h1E8FEA;
  c_a12[19] = 24'h197A49;
  c_a12[20] = 24'h15543B;
  c_a12[21] = 24'h11FEBA;
  c_a12[22] = 24'h0F61AE;
  c_a12[23] = 24'h0D6ACB;
  c_a12[24] = 24'h0C0CA7;
  c_a12[25] = 24'h0B3E1D;
  c_a12[26] = 24'h0AF9D9;
  c_a12[27] = 24'h0B3E1D;
  c_a12[28] = 24'h0C0CA7;
  c_a12[29] = 24'h0D6ACB;
  c_a12[30] = 24'h0F61AE;
  c_a12[31] = 24'h11FEBA;
  c_a12[32] = 24'h15543B;
  c_a12[33] = 24'h197A49;
  c_a12[34] = 24'h1E8FEA;
  c_a12[35] = 24'h3DAC66;
  c_a12[36] = 24'h3B6E74;
  c_a12[37] = 24'h373067;
  c_a12[38] = 24'h352ED0;
  c_a12[39] = 24'h333FE8;
  c_a12[40] = 24'h316303;
  c_a12[41] = 24'h2F977E;
  c_a12[42] = 24'h2DDCBA;
  c_a12[43] = 24'h2C3220;
  c_a12[44] = 24'h2A971F;
  c_a12[45] = 24'h290B2C;
  c_a12[46] = 24'h278DC4;
  c_a12[47] = 24'h261E66;
  c_a12[48] = 24'h24BC99;
  c_a12[49] = 24'h2367EA;
  c_a12[50] = 24'h221FE8;
  c_a12[51] = 24'h20E42B;
  c_a12[52] = 24'h1FB44C;
  c_a12[53] = 24'h1E8FEA;
  c_a12[54] = 24'h197A49;
  c_a12[55] = 24'h15543B;
  c_a12[56] = 24'h11FEBA;
  c_a12[57] = 24'h0F61AE;
  c_a12[58] = 24'h0D6ACB;
  c_a12[59] = 24'h0C0CA7;
  c_a12[60] = 24'h0B3E1D;
  c_a12[61] = 24'h0AF9D9;
  c_a12[62] = 24'h0B3E1D;
  c_a12[63] = 24'h0C0CA7;
  c_a12[64] = 24'h0D6ACB;
  c_a12[65] = 24'h0F61AE;
  c_a12[66] = 24'h11FEBA;
  c_a12[67] = 24'h15543B;
  c_a12[68] = 24'h197A49;
  c_a12[69] = 24'h1E8FEA;
  c_a12[70] = 24'h3DAC66;
  c_a12[71] = 24'h3B6E74;
  c_a12[72] = 24'h373067;
  c_a12[73] = 24'h352ED0;
  c_a12[74] = 24'h333FE8;
  c_a12[75] = 24'h316303;
  c_a12[76] = 24'h2F977E;
  c_a12[77] = 24'h2DDCBA;
  c_a12[78] = 24'h2C3220;
  c_a12[79] = 24'h2A971F;
  c_a12[80] = 24'h290B2C;
  c_a12[81] = 24'h278DC4;
  c_a12[82] = 24'h261E66;
  c_a12[83] = 24'h24BC99;
  c_a12[84] = 24'h2367EA;
  c_a12[85] = 24'h221FE8;
  c_a12[86] = 24'h20E42B;
  c_a12[87] = 24'h1FB44C;
  c_a12[88] = 24'h1E8FEA;
  c_a12[89] = 24'h197A49;
  c_a12[90] = 24'h15543B;
  c_a12[91] = 24'h11FEBA;
  c_a12[92] = 24'h0F61AE;
  c_a12[93] = 24'h0D6ACB;
  c_a12[94] = 24'h0C0CA7;
  c_a12[95] = 24'h0B3E1D;
  c_a12[96] = 24'h0AF9D9;
  c_a12[97] = 24'h0B3E1D;
  c_a12[98] = 24'h0C0CA7;
  c_a12[99] = 24'h0D6ACB;
  c_a12[100] = 24'h0F61AE;
  c_a12[101] = 24'h11FEBA;
  c_a12[102] = 24'h15543B;
  c_a12[103] = 24'h197A49;
  c_a12[104] = 24'h1E8FEA;

endfunction: setup_coefficients

task body;
  c_setup.rm = rm;
  setup_coefficients();

  cfg.mode = LP;
  for(int i = 0; i < 35; i++) begin
    c_setup.a11 = c_a11[i];
    c_setup.a12 = c_a12[i];
    c_setup.b10 = c_b10[i];
    c_setup.b11 = c_b11[i];
    c_setup.b12 = c_b12[i];
    c_setup.start(apb);
    `uvm_info("biquad_test::body", "Starting frequency sweep for new Low Pass filter configuration", UVM_LOW)
    f_sweep.start(signal);
  end

  cfg.mode = HP;
  for(int i = 35; i < 70; i++) begin
    c_setup.a11 = c_a11[i];
    c_setup.a12 = c_a12[i];
    c_setup.b10 = c_b10[i];
    c_setup.b11 = c_b11[i];
    c_setup.b12 = c_b12[i];
    c_setup.start(apb);
    `uvm_info("biquad_test::body", "Starting frequency sweep for new High Pass filter configuration", UVM_LOW)
    f_sweep.start(signal);
  end

  cfg.mode = BP;
  for(int i = 70; i < 105; i++) begin
    c_setup.a11 = c_a11[i];
    c_setup.a12 = c_a12[i];
    c_setup.b10 = c_b10[i];
    c_setup.b11 = c_b11[i];
    c_setup.b12 = c_b12[i];
    c_setup.start(apb);
    `uvm_info("biquad_test::body", "Starting frequency sweep for new Band Pass filter configuration", UVM_LOW)
    f_sweep.start(signal);
  end

endtask: body

endclass: biquad_vseq
