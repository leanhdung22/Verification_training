//
//------------------------------------------------------------------------------
//   Copyright 2018 Mentor Graphics Corporation
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//------------------------------------------------------------------------------
//
//------------------------------------------------------------------------------
//   Copyright 2018 Mentor Graphics Corporation
//   All Rights Reserved Worldwide
//
//   Licensed under the Apache License, Version 2.0 (the
//   "License"); you may not use this file except in
//   compliance with the License.  You may obtain a copy of
//   the License at
//
//       http://www.apache.org/licenses/LICENSE-2.0
//
//   Unless required by applicable law or agreed to in
//   writing, software distributed under the License is
//   distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
//   CONDITIONS OF ANY KIND, either express or implied.  See
//   the License for the specific language governing
//   permissions and limitations under the License.
//----- -------------------------------------------------------------------------
module sfr_dut #(ADDR_WIDTH = 8,
                 DATA_WIDTH = 8)
               (input clk,
                input reset,
                input[ADDR_WIDTH-1:0] address,
                input[DATA_WIDTH-1:0] write_data,
                input we,
                input re,
                output logic[DATA_WIDTH-1:0] read_data);

logic[DATA_WIDTH-1:0] mem[65535:0];

always @(posedge clk) begin
  begin
    if(we == 1) begin
      mem[address] = write_data;
    end
  end
end

always @(address or re) begin
  read_data = mem[address];
end

endmodule
