-------------------------------------------------------------------------------
-- Title      : vhdl_fsm
-- Project    : 
-------------------------------------------------------------------------------
-- File       : vhdl_fsm.vhd
-- Author     : LE  <le@le-VirtualBox>
-- Company    : 
-- Created    : 2019-02-06
-- Last update: 2019-02-06
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: cfg cours de VHDL SEI-2A-Phelma
-------------------------------------------------------------------------------
-- Copyright (c) 2019 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2019-02-06  1.0      le	Created
-------------------------------------------------------------------------------

-- C-cth: generating template infomation
